--
-- DLX_PROG2.vhd
--
-- Programa para el DLX32p
-- Se ha insertado nop para evitar las dependencias. Esta es la diferencia con DLX_PROG.vhd
-- que es el que se ha utilizado para DLX32s monociclo.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.DLX_pack.all;

package DLX_prog2 is
  type ROM_TABLE is array (0 to 88) of ROM_WORD;

  constant ROM: ROM_TABLE := ROM_TABLE'(

-- PROGRAMA PRINCIPAL
								--	; vector 1
--	ROM_WORD'("00110100000000010000000000010100"),  	--0	ORI R1, R0, 20
--	ROM_WORD'("00110100000000100000000000000010"),  	--4	ORI R2, R0, 2
	ROM_WORD'("00000000000000000000000000000000"),		--8	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--12	NOP
--	ROM_WORD'("00000000001000100001100000000111"),  	--16	SRA R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--20	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--24	NOP
--	ROM_WORD'("10101100000000110000000000000000"),  	--28	SW 0(R0), R3
--	ROM_WORD'("00000000000000000000000000000000"),		--32	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--36	NOP

--6 PRUEBAS ADELANTAMIENTO EN EX	
	ROM_WORD'("00110100000000010000000000010100"),  	--0	ORI R1, R0, 20
	ROM_WORD'("00110100000000100000000000000010"),  	--4	ORI R2, R0, 2
	ROM_WORD'("00000000001000100001100000000111"),  	--16	SRA R3, R1, R2
	ROM_WORD'("10101100000000110000000000000000"),  	--28	SW 0(R0), R3
	ROM_WORD'("00000000000000000000000000000000"),		--32	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--36	NOP

--8 PRUEBAS ADELANTAMIENTO DE CARGA - ALMACENAMIENTO
--	ROM_WORD'("10001100000000010000000000000000"),  	--320	LW 0(R0), R1
--	ROM_WORD'("10101100000000010000000000000000"),  	--320	SW 0(R0), R1
--	ROM_WORD'("00000000000000000000000000000000"),		--28	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--32	NOP
--	ROM_WORD'("10001100000000010000000000000000"),  	--320	LW 0(R0), R1
--	ROM_WORD'("00000000000000000000000000000000"),		--56	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00110100001000010000000000000000"),  	--40	ORI R1, R1, 0

--10 PRUEBAS ADELANTAMIENTO DE SALTOS CONDICIONALES
--	ROM_WORD'("00110110101101010000000000000001"),  	--40	ORI R21, R21, 1
--	ROM_WORD'("00010010101000000000000000010000"),  	--312	BEQZ R21, +16
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("00110111111111110000000000011100"),  	--40	ORI R31, R31, 28
--	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
--	ROM_WORD'("01001011111000000000000000000000"),  	--340	JR R31


	ROM_WORD'("00110100000000010000000000000100"),  	--40	ORI R1, R0, 4
	ROM_WORD'("00110100000000100000000000000011"),  	--44	ORI R2, R0, 3
	ROM_WORD'("00000000000000000000000000000000"),		--48	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--52	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--56	NOP
	ROM_WORD'("00000000001000100001100000000100"),  	--60	SLL R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--64	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--68	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--72	NOP
	ROM_WORD'("10101100000000110000000000000001"),  	--76	SW 1(R0), R3

	ROM_WORD'("00110100000000010000000000011000"),  	--80	ORI R1, R0, 24
	ROM_WORD'("00110100000000100000000000000010"),  	--84	ORI R2, R0, 2
	ROM_WORD'("00000000000000000000000000000000"),		--88	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--92	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--96	NOP
	ROM_WORD'("00000000001000100001100000000110"),  	--100	SRL R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--104	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--108	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--112	NOP
	ROM_WORD'("10101100000000110000000000000010"),  	--116	SW 2(R0), R3

								--	; vector 2
	ROM_WORD'("00110100000000010000000000000100"),  	--120	ORI R1, R0, 4
	ROM_WORD'("00110100000000100000000000001000"),  	--124	ORI R2, R0, 8
	ROM_WORD'("00000000000000000000000000000000"),		--128	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--132	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--136	NOP
	ROM_WORD'("00000000001000100001100000100101"),  	--140	OR R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--144	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--148	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--152	NOP
	ROM_WORD'("10101100000000110000000000000011"),  	--156	SW 3(R0), R3

	ROM_WORD'("00110100000000010000000000011100"),  	--160	ORI R1, R0, 28
	ROM_WORD'("00110100000000100000000000000011"),  	--164	ORI R2, R0, 3
	ROM_WORD'("00000000000000000000000000000000"),		--168	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--172	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--176	NOP
	ROM_WORD'("00000000001000100001100000100010"),  	--180	SUB R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--184	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--188	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--192	NOP
	ROM_WORD'("10101100000000110000000000000100"),  	--196	SW 4(R0), R3

	ROM_WORD'("00110100000000010000000000011000"),  	--200	ORI R1, R0, 24
	ROM_WORD'("00110100000000100000000000001000"),  	--204	ORI R2, R0, 8
	ROM_WORD'("00000000000000000000000000000000"),		--208	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--212	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--216	NOP
	ROM_WORD'("00000000001000100001100000100100"),  	--220	AND R3, R1, R2
	ROM_WORD'("00000000000000000000000000000000"),		--224	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--228	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--232	NOP
	ROM_WORD'("10101100000000110000000000000101"),  	--236	SW 5(R0), R3

								--	; llamadas al procedimiento
	ROM_WORD'("00001100000000000000000000110100"),  	--240	JAL SUMA_VECTOR ;(240 + 4 + 52 = 296)
	ROM_WORD'("00110100000111100000000000000000"),  	--244	ORI R30, R0, 0
	ROM_WORD'("00000000000111010000100000100000"),  	--248	ADD R1, R0, R29

	ROM_WORD'("00001100000000000000000000101000"),  	--252	JAL SUMA_VECTOR ;(252 + 4 + 40 = 296)
	ROM_WORD'("00110100000111100000000000000011"),  	--256	ORI R30, R0, 3
	ROM_WORD'("00000000000111010001000000100000"),  	--260	ADD R2, R0, R29
	ROM_WORD'("00000000000000000000000000000000"),		--264	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--268	NOP
	ROM_WORD'("00000000000000000000000000000000"),		--272	NOP

								--	; comparaci�n final
	ROM_WORD'("00000000001000100001100000101010"),  	--276	SLT R3, R1, R2

								--	; llamada al sistema, por ejemplo, escribir en pantalla el resultado
	ROM_WORD'("01000100000000000000000101011100"),  	--280	TRAP PANTALLA ;(348)
	ROM_WORD'("00000000000000000000000000000000"),		--284	NOP

								--	; finaliza la ejecuci�n del programa
	ROM_WORD'("01000100000000000000000000000000"),  	--288	TRAP 0
	ROM_WORD'("00000000000000000000000000000000"),		--292	NOP

-- FIN PROGRAMA PRINCIPAL

-- FUNCION SUMA_VECTOR

								--SUMA_VECTOR: ;(296) implemantaci�n del procedimiento 
								--	; inicializamos las variables locales
	ROM_WORD'("00110100000101010000000000000011"),  	--296	ORI R21, R0, 3 ; contador de iteraciones
	ROM_WORD'("00110100000101100000000000000001"),  	--300	ORI R22, R0, 1 ; decremento/incremento unidad
	ROM_WORD'("00110100000111010000000000000000"),  	--304	ORI R29, R0, 0 ; inicializaci�n del acumulado
	
								--LOOP: ;(308)
	ROM_WORD'("00000000000000000000000000000000"),		--308	NOP
	ROM_WORD'("00010010101000000000000000011000"),  	--312	BEQZ R21, END_LOOP ;(312 + 4 + 24 = 340)
	ROM_WORD'("00000000000000000000000000000000"),		--316	NOP
	ROM_WORD'("10001111110101110000000000000000"),  	--320	LW R23, 0(R30)
	ROM_WORD'("00000010101101101010100000100010"),  	--324	SUB R21, R21, R22
	ROM_WORD'("00000011110101101111000000100000"),  	--328	ADD R30, R30, R22
	ROM_WORD'("00001011111111111111111111100100"),  	--332	J LOOP ;(332 + 4 + (-28) = 308)
	ROM_WORD'("00000011101101111110100000100000"),  	--336	ADD R29, R29, R23
	
								--END_LOOP: ;(340) retornamos del procedimiento
	ROM_WORD'("01001011111000000000000000000000"),  	--340	JR R31	
	ROM_WORD'("00000000000000000000000000000000"),		--344	NOP
	
-- FIN FUNCION SUMA_VECTOR

-- LLAMADA AL SISTEMA
								--PANTALLA: ;(348) suponemos que ejecuta un syscall que escribe algo en pantalla
	ROM_WORD'("01000000000000000000000000000000"),  	--348	RFE			
	ROM_WORD'("00000000000000000000000000000000")		--352	NOP

-- FIN LLAMADA AL SISTEMA
      );

end DLX_prog2;


